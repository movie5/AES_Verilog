`timescale 1ns / 1ps

module GF_Multiplier(
    input [7:0] in1,
    input [7:0] in2,
    output [7:0] out
    );
    
//Modulo polynomials    
localparam modulo = 9'b100011011;

/***********************************



************************************/
endmodule
