`timescale 1ns / 1ps


module round_final(
    input [127:0] in
    );
    
    
endmodule
