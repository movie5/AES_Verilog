`timescale 1ns / 10ps

module ShiftRows_tb;

reg [127:0] in;
wire [127:0] out;

initial begin
    in = 128'hEA835CF00445332D655D98AD8596B0C5;
end

ShiftRows SR_1(in, out);

endmodule